library ieee;
  use ieee.std_logic_1164.all;

------------------------------------------------------------
-- Entity declaration for testbench
------------------------------------------------------------

entity top is
-- Entity of testbench is always empty
end entity top;

------------------------------------------------------------
-- Architecture body for testbench
------------------------------------------------------------

architecture testbench of top is

end architecture testbench;